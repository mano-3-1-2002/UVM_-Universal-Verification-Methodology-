`define DSIZE 8
`define ASIZE 4
